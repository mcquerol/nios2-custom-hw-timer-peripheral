
module customTimerPeripheral_tb();
